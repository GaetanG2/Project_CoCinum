
library ieee;
use ieee.std_logic_1164.all;

use work.Virgule_pkg.all;

entity UserInputs is
    generic(
        -- Declarations
    );
    port(
        -- Declarations
    );
end UserInputs;

architecture Behavioral of UserInputs is
    -- Declarations
begin
    -- Concurrent statements
end Behavioral;
