
library ieee;
use ieee.std_logic_1164.all;

use work.Virgule_pkg.all;

entity UserOutputs is
    generic(
        -- Declarations
    );
    port(
        -- Declarations
    );
end UserOutputs;

architecture Behavioral of UserOutputs is
    -- Declarations
begin
    -- Concurrent statements
end Behavioral;
